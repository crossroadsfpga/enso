// dc_fifo_convert_data_format_adapter_0.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module data_adapter (
		input  wire         clk,               //   clk.clk
		input  wire         reset_n,           // reset.reset_n
		input  wire [511:0] in_data,           //    in.data
		input  wire         in_valid,          //      .valid
		output wire         in_ready,          //      .ready
		input  wire         in_startofpacket,  //      .startofpacket
		input  wire         in_endofpacket,    //      .endofpacket
		input  wire [5:0]   in_empty,          //      .empty
		output wire [255:0] out_data,          //   out.data
		output wire         out_valid,         //      .valid
		input  wire         out_ready,         //      .ready
		output wire         out_startofpacket, //      .startofpacket
		output wire         out_endofpacket,   //      .endofpacket
		output wire [4:0]   out_empty          //      .empty
	);

	data_adapter_core data_adapter_core_0 (
		.clk               (clk),               //   input,    width = 1,   clk.clk
		.reset_n           (reset_n),           //   input,    width = 1, reset.reset_n
		.in_data           (in_data),           //   input,  width = 512,    in.data
		.in_valid          (in_valid),          //   input,    width = 1,      .valid
		.in_ready          (in_ready),          //  output,    width = 1,      .ready
		.in_startofpacket  (in_startofpacket),  //   input,    width = 1,      .startofpacket
		.in_endofpacket    (in_endofpacket),    //   input,    width = 1,      .endofpacket
		.in_empty          (in_empty),          //   input,    width = 6,      .empty
		.out_data          (out_data),          //  output,  width = 256,   out.data
		.out_valid         (out_valid),         //  output,    width = 1,      .valid
		.out_ready         (out_ready),         //   input,    width = 1,      .ready
		.out_startofpacket (out_startofpacket), //  output,    width = 1,      .startofpacket
		.out_endofpacket   (out_endofpacket),   //  output,    width = 1,      .endofpacket
		.out_empty         (out_empty)          //  output,    width = 5,      .empty
	);

endmodule
