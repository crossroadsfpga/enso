// dsp.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module dsp (
		input  wire [17:0] ay,      //      ay.ay
		input  wire [17:0] by,      //      by.by
		input  wire [17:0] ax,      //      ax.ax
		input  wire [17:0] bx,      //      bx.bx
		output wire [36:0] resulta, // resulta.resulta
		input  wire        clk0,    //    clk0.clk
		input  wire        clk1,    //    clk1.clk
		input  wire        clk2,    //    clk2.clk
		input  wire [2:0]  ena      //     ena.ena
	);

	dsp_altera_s10_native_fixed_point_dsp_181_5337kly s10_native_fixed_point_dsp_0 (
		.ay      (ay),      //   input,  width = 18,      ay.ay
		.by      (by),      //   input,  width = 18,      by.by
		.ax      (ax),      //   input,  width = 18,      ax.ax
		.bx      (bx),      //   input,  width = 18,      bx.bx
		.resulta (resulta), //  output,  width = 37, resulta.resulta
		.clk0    (clk0),    //   input,   width = 1,    clk0.clk
		.clk1    (clk1),    //   input,   width = 1,    clk1.clk
		.clk2    (clk2),    //   input,   width = 1,    clk2.clk
		.ena     (ena)      //   input,   width = 3,     ena.ena
	);

endmodule
